FOOTBALL_API_KEY ="dd82933e09e4052c68aafecf1feb4634"
SNOWFLAKE_ACCOUNT="RY83976.ap-southeast-1"
SNOWFLAKE_USER="LASTTIME1"
SNOWFLAKE_PASSWORD="Maxttime1@tawan"
SNOWFLAKE_WAREHOUSE="COMPUTE_WH"
SNOWFLAKE_DATABASE="FOOTBALL_CAPSTONE"
SNOWFLAKE_SCHEMA="RAW"
SNOWFLAKE_ROLE="ACCOUNTADMIN"


Github = "https://github.com/tawanwetaya-debug/Capstone---Football.git"

