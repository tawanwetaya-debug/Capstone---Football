FOOTBALL_API_KEY ="dd82933e09e4052c68aafecf1feb4634"
SNOWFLAKE_ACCOUNT="WOIQSGO-AJ77687"
SNOWFLAKE_USER="LASTTIME2"
SNOWFLAKE_PASSWORD="Maxttime1@tawan"
SNOWFLAKE_WAREHOUSE="COMPUTE_WH"
SNOWFLAKE_DATABASE="FOOTBALL_CAPSTONE"
SNOWFLAKE_SCHEMA="RAW"
SNOWFLAKE_ROLE="ACCOUNTADMIN"


Github = "https://github.com/tawanwetaya-debug/Capstone---Football.git"

